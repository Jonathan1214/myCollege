module MEM ;

endmodule

module SC;

endmodule

module Xbar;

endmodule
