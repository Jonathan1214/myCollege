module IS;
    MEM mem1;
    SC sc1;
    Xbar xbar1;
endmodule