module FA;
endmodule