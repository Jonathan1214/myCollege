module Top;
    IS is1;
endmodule